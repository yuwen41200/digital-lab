/**
 * Rotary Dial Controller
 * Copyright Notice: This code was written by the TAs of this course.
 */

module rotary_ctrl(
		input rst,
		input clk,
		input rot_a,
		input rot_b,
		output [7:0] led
	);

endmodule
